/*************************************************************************
 > Copyright (C) 2021 Sangfor Ltd. All rights reserved.
 > File Name   : wshb_bfm_pkg.sv
 > Author      : bhyou
 > Mail        : bhyou@foxmail.com 
 > Created Time: Sun 26 Dec 2021 02:04:02 PM CST
 ************************************************************************/
 
package wshb_bfn_pkg;


    
endpackage